`timescale 1ns / 1ps

module tb_ultrasonic();
    reg clk;
    reg reset;
    reg echo;
    wire trigger;
    wire [8:0] distance;

    ultrasonic_sensor u_ultra_tb(
        .clk(clk),
        .reset(reset),
        .echo(echo),
        .trigger(trigger),
        .distance(distance)
    );

    initial begin
        clk = 0;
        reset = 1;
        echo = 0;
    end


    always #5 clk = ~clk;

    initial begin
        #10 reset = 0;
        #10 wait(trigger); // wait 1    // when state = S_T_HIGH_10, 16us trigger transmit / wait trigger pedge
             wait(!trigger); // wiat 0  // when finish 16us trigger transmit / wait trigger nedge / 
        #20000; // wait 20us
        echo = 1; #800000; // wait // echo 800us => 13 cm
        echo = 0;
        #10000; $stop;
    end


endmodule
